`timescale 1ns/1ps
// -----------------------------------------------------------------------------
// ISO‑16 True Delivery Loop — Reference RTL (informative)
// -----------------------------------------------------------------------------
// This module is an informative, non‑normative reference implementation of the
// ISO‑16 True Delivery Loop state machine. It is intended as a behavioral and
// timing oracle for vendors and auditors.
//
// Normative behavior is defined by the written specification, conformance
// vectors, and Golden Waveform templates. If a discrepancy is found, the
// written specification prevails.
// -----------------------------------------------------------------------------

module iso16_true_delivery #(
    parameter integer NUM_PLUGINS   = 4,
    parameter integer WARP_WIDTH    = 16,   // Q16.16 or similar
    parameter integer ERROR_WIDTH   = 32,
    parameter integer LATTICE_SIZE  = 16    // 4x4 lattice flattened
)(
    input  wire                     clk,
    input  wire                     rst_n,
    input  wire                     start,
    input  wire [15:0]              vector_id,
    input  wire [ERROR_WIDTH-1:0]   epsilon,

    // Plugin interface (flattened buses for Verilog‑2001 compatibility)
    input  wire [NUM_PLUGINS-1:0]                       plugin_valid,
    input  wire [NUM_PLUGINS*WARP_WIDTH-1:0]           plugin_warp_x,
    input  wire [NUM_PLUGINS*WARP_WIDTH-1:0]           plugin_warp_y,
    input  wire [NUM_PLUGINS*WARP_WIDTH-1:0]           plugin_warp_z,
    input  wire [NUM_PLUGINS*ERROR_WIDTH-1:0]          plugin_error,

    // State machine visibility
    output reg  [2:0]               state,

    // Accumulators
    output reg  [WARP_WIDTH-1:0]    warp_sum_x,
    output reg  [WARP_WIDTH-1:0]    warp_sum_y,
    output reg  [WARP_WIDTH-1:0]    warp_sum_z,
    output reg  [ERROR_WIDTH-1:0]   error_sum,

    // Check results
    output reg                      symmetry_ok,
    output reg                      error_ok,
    output reg                      true_delivery,

    // Seal boundary
    output reg                      seal_start,
    output reg                      seal_ready,
    output reg  [255:0]             seal
);

    // -------------------------------------------------------------------------
    // State machine encoding
    // -------------------------------------------------------------------------
    localparam [2:0]
        ST_IDLE       = 3'd0,
        ST_COLLECT    = 3'd1,
        ST_ACCUMULATE = 3'd2,
        ST_APPLY      = 3'd3,
        ST_CHECK      = 3'd4,
        ST_SEAL       = 3'd5,
        ST_DONE       = 3'd6;

    reg [2:0] state_next;

    // -------------------------------------------------------------------------
    // Canonical lattice (informative ROM)
    // 4x4 lattice flattened to 16 entries. Values are placeholders; in a
    // complete reference, these would be the canonical Q16.16 coordinates.
    // -------------------------------------------------------------------------
    reg [WARP_WIDTH-1:0] canonical_lattice_x [0:LATTICE_SIZE-1];
    reg [WARP_WIDTH-1:0] canonical_lattice_y [0:LATTICE_SIZE-1];
    reg [WARP_WIDTH-1:0] canonical_lattice_z [0:LATTICE_SIZE-1];

    initial begin : init_lattice
        integer i;
        for (i = 0; i < LATTICE_SIZE; i = i + 1) begin
            canonical_lattice_x[i] = {WARP_WIDTH{1'b0}};
            canonical_lattice_y[i] = {WARP_WIDTH{1'b0}};
            canonical_lattice_z[i] = {WARP_WIDTH{1'b0}};
        end
        // If you have specific canonical coordinates, assign them here.
    end

    // Warped lattice
    reg [WARP_WIDTH-1:0] phase_warped_x [0:LATTICE_SIZE-1];
    reg [WARP_WIDTH-1:0] phase_warped_y [0:LATTICE_SIZE-1];
    reg [WARP_WIDTH-1:0] phase_warped_z [0:LATTICE_SIZE-1];

    // -------------------------------------------------------------------------
    // Helper: extract plugin fields from flattened buses
    // -------------------------------------------------------------------------
    function [WARP_WIDTH-1:0] get_warp_x;
        input integer idx;
        begin
            get_warp_x = plugin_warp_x[idx*WARP_WIDTH +: WARP_WIDTH];
        end
    endfunction

    function [WARP_WIDTH-1:0] get_warp_y;
        input integer idx;
        begin
            get_warp_y = plugin_warp_y[idx*WARP_WIDTH +: WARP_WIDTH];
        end
    endfunction

    function [WARP_WIDTH-1:0] get_warp_z;
        input integer idx;
        begin
            get_warp_z = plugin_warp_z[idx*WARP_WIDTH +: WARP_WIDTH];
        end
    endfunction

    function [ERROR_WIDTH-1:0] get_error;
        input integer idx;
        begin
            get_error = plugin_error[idx*ERROR_WIDTH +: ERROR_WIDTH];
        end
    endfunction

    // -------------------------------------------------------------------------
    // Accumulation (COMB) — warp_sum and error_sum
    // -------------------------------------------------------------------------
    reg [WARP_WIDTH-1:0]    warp_sum_x_next;
    reg [WARP_WIDTH-1:0]    warp_sum_y_next;
    reg [WARP_WIDTH-1:0]    warp_sum_z_next;
    reg [ERROR_WIDTH-1:0]   error_sum_next;

    integer i;

    always @* begin
        warp_sum_x_next = {WARP_WIDTH{1'b0}};
        warp_sum_y_next = {WARP_WIDTH{1'b0}};
        warp_sum_z_next = {WARP_WIDTH{1'b0}};
        error_sum_next  = {ERROR_WIDTH{1'b0}};

        if (state == ST_ACCUMULATE) begin
            for (i = 0; i < NUM_PLUGINS; i = i + 1) begin
                if (plugin_valid[i]) begin
                    warp_sum_x_next = warp_sum_x_next + get_warp_x(i);
                    warp_sum_y_next = warp_sum_y_next + get_warp_y(i);
                    warp_sum_z_next = warp_sum_z_next + get_warp_z(i);
                    error_sum_next  = error_sum_next  + get_error(i);
                end
            end
        end
    end

    // -------------------------------------------------------------------------
    // APPLY: warp lattice (SEQ)
    // -------------------------------------------------------------------------
    integer j;

    // -------------------------------------------------------------------------
    // Symmetry check (COMB)
    // For simplicity, compare symmetric pairs (0,15), (1,14), ..., (7,8).
    // In a full reference, this should match the exact symmetry definition.
    // -------------------------------------------------------------------------
    reg symmetry_ok_next;

    always @* begin
        symmetry_ok_next = 1'b1;
        if (state == ST_CHECK) begin
            for (j = 0; j < LATTICE_SIZE/2; j = j + 1) begin
                if (phase_warped_x[j] != phase_warped_x[LATTICE_SIZE-1-j]) symmetry_ok_next = 1'b0;
                if (phase_warped_y[j] != phase_warped_y[LATTICE_SIZE-1-j]) symmetry_ok_next = 1'b0;
                if (phase_warped_z[j] != phase_warped_z[LATTICE_SIZE-1-j]) symmetry_ok_next = 1'b0;
            end
        end
    end

    // -------------------------------------------------------------------------
    // Error check (COMB)
    // -------------------------------------------------------------------------
    reg error_ok_next;

    always @* begin
        error_ok_next = 1'b0;
        if (state == ST_CHECK) begin
            error_ok_next = (error_sum <= epsilon);
        end
    end

    // -------------------------------------------------------------------------
    // True delivery (COMB)
    // -------------------------------------------------------------------------
    reg true_delivery_next;

    always @* begin
        true_delivery_next = 1'b0;
        if (state == ST_CHECK) begin
            true_delivery_next = symmetry_ok_next & error_ok_next;
        end
    end

    // -------------------------------------------------------------------------
    // Seal engine interface (informative)
    // This module assumes an external SHA3‑256 core with a simple handshake.
//  The core is not defined here; this module focuses on seal boundary timing.
// -------------------------------------------------------------------------
    reg         seal_start_next;
    reg         seal_ready_next;
    reg [255:0] seal_next;

    // Simple illustrative behavior:
    // - On ST_SEAL entry, pulse seal_start for one cycle.
    // - After a fixed latency (e.g., 8 cycles), assert seal_ready and
    //   present a deterministic "digest" derived from internal state.
    //
    // In a complete reference, this would drive a real SHA3‑256 core and
    // serialize the canonical fields as defined in the spec.

    localparam integer SEAL_LATENCY = 8;
    reg [3:0] seal_counter;

    always @* begin
        seal_start_next = 1'b0;
        seal_ready_next = seal_ready;
        seal_next       = seal;

        if (state == ST_SEAL) begin
            if (seal_counter == 0) begin
                // First cycle in SEAL: start seal
                seal_start_next = 1'b1;
            end
        end
    end

    // -------------------------------------------------------------------------
    // State machine + sequential logic
    // -------------------------------------------------------------------------
    always @* begin
        state_next = state;
        case (state)
            ST_IDLE: begin
                if (start)
                    state_next = ST_COLLECT;
            end

            ST_COLLECT: begin
                // Plugins present stable data during this window.
                state_next = ST_ACCUMULATE;
            end

            ST_ACCUMULATE: begin
                state_next = ST_APPLY;
            end

            ST_APPLY: begin
                state_next = ST_CHECK;
            end

            ST_CHECK: begin
                state_next = ST_SEAL;
            end

            ST_SEAL: begin
                if (seal_counter == SEAL_LATENCY)
                    state_next = ST_DONE;
            end

            ST_DONE: begin
                // One‑shot; return to IDLE when start is deasserted and reasserted.
                if (!start)
                    state_next = ST_IDLE;
            end

            default: state_next = ST_IDLE;
        endcase
    end

    // Sequential block
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state         <= ST_IDLE;
            warp_sum_x    <= {WARP_WIDTH{1'b0}};
            warp_sum_y    <= {WARP_WIDTH{1'b0}};
            warp_sum_z    <= {WARP_WIDTH{1'b0}};
            error_sum     <= {ERROR_WIDTH{1'b0}};
            symmetry_ok   <= 1'b0;
            error_ok      <= 1'b0;
            true_delivery <= 1'b0;
            seal_start    <= 1'b0;
            seal_ready    <= 1'b0;
            seal          <= 256'h0;
            seal_counter  <= 4'd0;

            for (j = 0; j < LATTICE_SIZE; j = j + 1) begin
                phase_warped_x[j] <= {WARP_WIDTH{1'b0}};
                phase_warped_y[j] <= {WARP_WIDTH{1'b0}};
                phase_warped_z[j] <= {WARP_WIDTH{1'b0}};
            end
        end else begin
            state <= state_next;

            // Accumulators latch at end of ACCUMULATE
            if (state == ST_ACCUMULATE) begin
                warp_sum_x <= warp_sum_x_next;
                warp_sum_y <= warp_sum_y_next;
                warp_sum_z <= warp_sum_z_next;
                error_sum  <= error_sum_next;
            end

            // APPLY: warp lattice
            if (state == ST_APPLY) begin
                for (j = 0; j < LATTICE_SIZE; j = j + 1) begin
                    phase_warped_x[j] <= canonical_lattice_x[j] + warp_sum_x_next;
                    phase_warped_y[j] <= canonical_lattice_y[j] + warp_sum_y_next;
                    phase_warped_z[j] <= canonical_lattice_z[j] + warp_sum_z_next;
                end
            end

            // CHECK: latch results
            if (state == ST_CHECK) begin
                symmetry_ok   <= symmetry_ok_next;
                error_ok      <= error_ok_next;
                true_delivery <= true_delivery_next;
            end

            // SEAL timing
            if (state == ST_SEAL) begin
                seal_start <= seal_start_next;

                if (seal_counter < SEAL_LATENCY)
                    seal_counter <= seal_counter + 1'b1;

                if (seal_counter == SEAL_LATENCY) begin
                    seal_ready <= 1'b1;
                    // Deterministic placeholder digest derived from internal state.
                    // In a full reference, this would be the SHA3‑256 of the
                    // canonical serialization.
                    seal <= {
                        vector_id,
                        warp_sum_x,
                        warp_sum_y,
                        warp_sum_z,
                        error_sum[31:0],
                        16'h0000,
                        8'h00,
                        symmetry_ok,
                        error_ok,
                        true_delivery,
                        215'd0
                    };
                end
            end else begin
                seal_start   <= 1'b0;
                seal_ready   <= 1'b0;
                seal_counter <= 4'd0;
            end
        end
    end

endmodule
